--
-- VHDL Architecture Cursor_test.CursorMaster_tester.test
--
-- Created:
--          by - Arnaud.UNKNOWN (DESKTOP-4F3HILT)
--          at - 14:20:09 06.12.2021
--
-- using Mentor Graphics HDL Designer(TM) 2019.2 (Build 5)
--
ARCHITECTURE test OF CursorMaster_tester IS
BEGIN
END ARCHITECTURE test;

